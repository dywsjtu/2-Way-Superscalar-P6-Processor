`ifndef __FU_MULT_V__
`define __FU_MULT_V__

`timescale 1ns/100ps

module fu_mult(
	input                           clock,               // system clock
	input                           reset,               // system reset
	input							valid,
    input	ID_RS_PACKET			id_fu,
	input   RS_FU_PACKET            rs_fu,

    output  FU_RS_PACKET            fu_rs,
	output							fu_result_valid
);
	logic 	[`XLEN-1:0] 			opa_mux_out, opb_mux_out;
	logic	[`XLEN-1:0]				alu_result;
    logic                           alu_result_valid;
	ID_RS_PACKET					working_id_fu;
	RS_FU_PACKET					working_rs_fu;

	// Pass-throughs
	assign fu_rs.NPC            = working_id_fu.NPC;
	assign fu_rs.rs2_value      = working_rs_fu.rs_value[1];
	assign fu_rs.rd_mem         = working_id_fu.rd_mem;
	assign fu_rs.wr_mem         = working_id_fu.wr_mem;
	assign fu_rs.dest_reg_idx   = working_id_fu.dest_reg_idx;
	assign fu_rs.halt           = working_id_fu.halt;
	assign fu_rs.illegal        = working_id_fu.illegal;
	assign fu_rs.csr_op         = working_id_fu.csr_op;
	assign fu_rs.mem_size       = working_id_fu.inst.r.funct3;
	assign fu_result_valid		= ~working_rs_fu.selected &&
								  working_id_fu.valid && working_rs_fu.rs_value_valid && 
								  alu_result_valid;
	
	//
	// ALU opA mux
	//
	assign opa_mux_out = working_rs_fu.rs_value[0];

	//
	// ALU opB mux
	//
	assign opb_mux_out = working_rs_fu.rs_value[1];

	//
	// instantiate the ALU
	//
	mlu mlu_0 (// Inputs
		.clock(clock),
		.reset(reset),

		.refresh(working_rs_fu.squash || working_rs_fu.selected),
		.val_valid(working_rs_fu.rs_value_valid),
		.opa(opa_mux_out),
		.opb(opb_mux_out),
		.func(working_id_fu.alu_func),

		// Output
		.valid(alu_result_valid),
		.result(alu_result)
	);

	 // ultimate "take branch" signal:
	 //	unconditional, or conditional and the condition is true
	assign fu_rs.take_branch = 1'b0;
	assign fu_rs.alu_result	 = alu_result;

	// synopsys sync_set_reset "reset"
	always_ff @(posedge clock) begin
		if (reset || rs_fu.squash) begin
			working_id_fu				<=	`SD	0;
			working_rs_fu				<=	`SD	0;
		end else if (rs_fu.selected) begin
			if (valid && id_fu.valid && id_fu.dispatch_enable) begin
				working_id_fu			<=	`SD	id_fu;
				working_rs_fu.squash		<=	`SD	rs_fu.squash;
				working_rs_fu.selected		<=	`SD	1'b1;
				working_rs_fu.rs_value		<=	`SD rs_fu.rs_value;
				working_rs_fu.rs_value_valid<=	`SD rs_fu.rs_value_valid;
			end else begin
				working_id_fu			<=	`SD	0;
				working_rs_fu			<=	`SD	{	1'b0,
													1'b1,
													{`XLEN'b0, `XLEN'b0},
													1'b0	};
			end
		end else begin
			if (valid && id_fu.valid && id_fu.dispatch_enable && ~working_id_fu.valid) begin
				working_id_fu				<=	`SD	id_fu;
				working_rs_fu.squash		<=	`SD	rs_fu.squash;
				working_rs_fu.selected		<=	`SD	1'b1;
				working_rs_fu.rs_value		<=	`SD rs_fu.rs_value;
				working_rs_fu.rs_value_valid<=	`SD rs_fu.rs_value_valid;
			end else begin 
				if (working_id_fu.valid && rs_fu.rs_value_valid && ~working_rs_fu.rs_value_valid) begin
					// working_rs_fu			<=	`SD	rs_fu;
					working_rs_fu.squash		<=	`SD	rs_fu.squash;
					working_rs_fu.selected		<=	`SD	1'b1;
					working_rs_fu.rs_value		<=	`SD rs_fu.rs_value;
					working_rs_fu.rs_value_valid<=	`SD rs_fu.rs_value_valid;
				end else if (working_rs_fu.selected) begin
					working_rs_fu.selected	<=	`SD	1'b0;
				end
			end
		end
	end

endmodule // module fu_mult
`endif // __FU_MULT_V__
